-- Adder 

LIBRARY sxlib_ModelSim;

ENTITY  alu IS
  PORT (
		a 	: in bit_vector(3 downto 0);
		b 	: in bit_vector(3 downto 0);
		s	: out bit_vector(3 downto 0);
                vdd     : in bit;
                vss     : in bit
    );
END  alu;

-- Architecture Declaration

ARCHITECTURE behaviour_data_flow OF  alu IS

-- carry

  SIGNAL carry : BIT_VECTOR(3 downto 0) ;

BEGIN

-- carru definition

carry(0) <= '0';
carry(3 downto 1) <= ( ( b(2 downto 0) and a(2 downto 0) ) or
                   ( a(2 downto 0) and carry(2 downto 0) ) or
		   ( carry(2 downto 0) and b(2 downto 0) ) ) ;

-- sum definition

s <= b xor a xor carry ;

END;


-- Architecture Declaration

ARCHITECTURE structural_view OF alu IS

  COMPONENT a2_x2
    port (
	  i0 : in BIT;        -- i0
	  i1 : in BIT;        -- i1
	  q : out BIT;        -- t
	  vdd : in BIT;       -- vdd
	  vss : in BIT        -- vss
    );
  END COMPONENT;

  COMPONENT o3_x2
    port (
    i0 : in BIT;        -- i0
    i1 : in BIT;        -- i1
    i2 : in BIT;        -- i2
    q  : out BIT;        -- f
    vdd : in BIT;       -- vdd
    vss : in BIT        -- vss
    );
  END COMPONENT;

  COMPONENT xr2_x1
PORT (
  i0	 : in  BIT;
  i1	 : in  BIT;
  q	 : out BIT;
  vdd	 : in  BIT;
  vss	 : in  BIT
);
  END COMPONENT;

-- carry signals	

  SIGNAL carry   : bit_vector (2 downto 0);
  signal carry_0 : bit_vector (2 downto 1);
  signal carry_1 : bit_vector (2 downto 1);
  signal carry_2 : bit_vector (2 downto 1);
  signal sum : bit_vector (3 downto 1);

BEGIN

-- instances

  carry_0_0  : a2_x2 port map(b(0), a(0), carry(0), vdd, vss);
  carry_0_1  : a2_x2 port map(b(1), a(1), carry_0(1), vdd, vss);
  carry_0_2  : a2_x2 port map(b(2), a(2), carry_0(2), vdd, vss);

  carry_1_1  : a2_x2 port map(b(1), carry(0), carry_1(1), vdd, vss);
  carry_1_2  : a2_x2 port map(b(2), carry(1), carry_1(2), vdd, vss);
  carry_2_1  : a2_x2 port map(a(1), carry(0), carry_2(1), vdd, vss);
  carry_2_2  : a2_x2 port map(a(2), carry(1), carry_2(2), vdd, vss);

  carry_out_1: o3_x2 port map(carry_0(1), carry_1(1), carry_2(1), carry(1), vdd, vss);
  carry_out_2: o3_x2 port map(carry_0(2), carry_1(2), carry_2(2), carry(2), vdd, vss);

  sum_0_0 : xr2_x1 port map(a(0), b(0), s(0), vdd, vss);
  sum_0_1 : xr2_x1 port map(a(1), b(1), sum(1), vdd, vss);
  sum_0_2 : xr2_x1 port map(a(2), b(2), sum(2), vdd, vss);
  sum_0_3 : xr2_x1 port map(a(3), b(3), sum(3), vdd, vss);

  sum_1_1 : xr2_x1 port map(sum(1), carry(0), s(1), vdd, vss);
  sum_1_2 : xr2_x1 port map(sum(2), carry(1), s(2), vdd, vss);
  sum_1_3 : xr2_x1 port map(sum(3), carry(2), s(3), vdd, vss);

end structural_view;
